`timescale 1ns / 1ps

// Generated ALU Module
// Style: STANDARD
// Bit width: 32
// Operations: ADD, SUB, AND, OR, XNOR, PASSB, XOR, ROL
// Flags: carry, zero, overflow, sign

module ALU_0455W32_4b0875b4(
    input  wire [3:0]  opcode,
    input  wire [31:0] input1,
    input  wire [31:0] input2,
    input  wire [4:0]       shiftValue,
    output wire [31:0] result
    ,output wire carryFlag
    ,output wire zeroFlag
    ,output wire overFlowFlag
    ,output wire signFlag
);

    // Operation codes
    localparam ADD = 4'd0;
    localparam SUB = 4'd1;
    localparam AND = 4'd2;
    localparam OR = 4'd3;
    localparam XNOR = 4'd4;
    localparam PASSB = 4'd5;
    localparam XOR = 4'd6;
    localparam ROL = 4'd7;

    // Internal signals
    wire [32:0] sum = (opcode == SUB) ? 
                             {1'b0, input1} - {1'b0, input2} : 
                             {1'b0, input1} + {1'b0, input2};

    // Combinational logic
    always @(*) begin
        case (opcode)
            ADD: begin
                result = input1 + input2;
                overflow = (input1[31] == input2[31]) && (result[31] != input1[31]);
            end
            SUB: begin
                result = input1 - input2;
                overflow = (input1[31] != input2[31]) && (result[31] != input1[31]);
            end
            AND: begin
                result = input1 & input2;
            end
            OR: begin
                result = input1 | input2;
            end
            XNOR: begin
                result = ~(input1 ^ input2);
            end
            PASSB: begin
                result = input2;
            end
            XOR: begin
                result = input1 ^ input2;
            end
            ROL: begin
                result = rol(input1, shiftValue);
            end
            default: result = 32'b0;
        endcase
        zeroFlag = (result == 32'b0);
        signFlag = result[31];
    end

endmodule