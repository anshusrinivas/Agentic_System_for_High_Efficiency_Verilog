`timescale 1ns / 1ps

// Generated ALU Module
// Style: OPTIMIZED
// Bit width: 32
// Operations: ADD, SUB, AND, OR, SLL, XOR, MUL, PASSB, NOR, SLT, ROL, SRA
// Flags: carry, zero, overflow, sign

module ALU_0277W32_b962a36b(
    input  wire [3:0]  opcode,
    input  wire [31:0] input1,
    input  wire [31:0] input2,
    input  wire [4:0]       shiftValue,
    output reg  [31:0] result
    ,output reg  carryFlag
    ,output reg  zeroFlag
    ,output reg  overFlowFlag
    ,output reg  signFlag
);

    // Operation codes
    localparam ADD = 4'd0;
    localparam SUB = 4'd1;
    localparam AND = 4'd2;
    localparam OR = 4'd3;
    localparam SLL = 4'd4;
    localparam XOR = 4'd5;
    localparam MUL = 4'd6;
    localparam PASSB = 4'd7;
    localparam NOR = 4'd8;
    localparam SLT = 4'd9;
    localparam ROL = 4'd10;
    localparam SRA = 4'd11;

    // Internal signals
    wire [32:0] sum = (opcode == SUB) ? 
                             {1'b0, input1} - {1'b0, input2} : 
                             {1'b0, input1} + {1'b0, input2};

    // Combinational logic
    always @(*) begin
        case (opcode)
            ADD: begin
                result = input1 + input2;
                overflow = (input1[31] == input2[31]) && (result[31] != input1[31]);
            end
            SUB: begin
                result = input1 - input2;
                overflow = (input1[31] != input2[31]) && (result[31] != input1[31]);
            end
            AND: begin
                result = input1 & input2;
            end
            OR: begin
                result = input1 | input2;
            end
            SLL: begin
                result = input1 << shiftValue;
            end
            XOR: begin
                result = input1 ^ input2;
            end
            MUL: begin
                result = input1 * input2;
            end
            PASSB: begin
                result = input2;
            end
            NOR: begin
                result = ~(input1 | input2);
            end
            SLT: begin
            end
            ROL: begin
                result = rol(input1, shiftValue);
            end
            SRA: begin
                result = $signed(input1) >>> shiftValue;
            end
            default: result = 32'b0;
        endcase
        zeroFlag = (result == 32'b0);
        signFlag = result[31];
    end

endmodule