`timescale 1ns / 1ps

// Generated ALU Module
// Style: STANDARD
// Bit width: 8
// Operations: ADD, SUB, AND, OR, PASSB, SRA, NAND, MAX
// Flags: carry

module ALU_1480W8_d18f8bcf(
    input  wire [3:0]  opcode,
    input  wire [7:0] input1,
    input  wire [7:0] input2,
    input  wire [4:0]       shiftValue,
    output wire [7:0] result
    ,output wire carryFlag
);

    // Operation codes
    localparam ADD = 4'd0;
    localparam SUB = 4'd1;
    localparam AND = 4'd2;
    localparam OR = 4'd3;
    localparam PASSB = 4'd4;
    localparam SRA = 4'd5;
    localparam NAND = 4'd6;
    localparam MAX = 4'd7;

    // Internal signals
    wire [8:0] sum = (opcode == SUB) ? 
                             {1'b0, input1} - {1'b0, input2} : 
                             {1'b0, input1} + {1'b0, input2};

    // Combinational logic
    always @(*) begin
        case (opcode)
            ADD: begin
                result = input1 + input2;
                
            end
            SUB: begin
                result = input1 - input2;
                
            end
            AND: begin
                result = input1 & input2;
            end
            OR: begin
                result = input1 | input2;
            end
            PASSB: begin
                result = input2;
            end
            SRA: begin
                result = $signed(input1) >>> shiftValue;
            end
            NAND: begin
                result = ~(input1 & input2);
            end
            MAX: begin
                result = (input1 > input2) ? input1 : input2;
            end
            default: result = 8'b0;
        endcase
    end

endmodule