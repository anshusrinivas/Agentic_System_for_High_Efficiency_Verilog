`timescale 1ns / 1ps

// Generated ALU Module
// Style: FUNCTION
// Bit width: 8
// Operations: ROL, ROR, MAX, MIN, ADD, SLL, SUB, XOR, XNOR, SRA
// Flags: carry, zero, overflow, sign

module ALU_0026W8_7ac7dc9f(
    input  wire [3:0]  opcode,
    input  wire [7:0] input1,
    input  wire [7:0] input2,
    input  wire [4:0]       shiftValue,
    output wire [7:0] result
    ,output wire carryFlag
    ,output wire zeroFlag
    ,output wire overFlowFlag
    ,output wire signFlag
);

    function [7:0] rol;
        input [7:0] a;
        input [4:0] sh;
        begin
            rol = (a << sh) | (a >> (8-sh));
        end
    endfunction

    function [7:0] ror;
        input [7:0] a;
        input [4:0] sh;
        begin
            ror = (a >> sh) | (a << (8-sh));
        end
    endfunction

    // Operation codes
    localparam ROL = 4'd0;
    localparam ROR = 4'd1;
    localparam MAX = 4'd2;
    localparam MIN = 4'd3;
    localparam ADD = 4'd4;
    localparam SLL = 4'd5;
    localparam SUB = 4'd6;
    localparam XOR = 4'd7;
    localparam XNOR = 4'd8;
    localparam SRA = 4'd9;

    // Internal signals
    wire [8:0] sum = (opcode == SUB) ? 
                             {1'b0, input1} - {1'b0, input2} : 
                             {1'b0, input1} + {1'b0, input2};

    // Combinational logic
    always @(*) begin
        case (opcode)
            ROL: begin
                result = rol(input1, shiftValue);
            end
            ROR: begin
                result = ror(input1, shiftValue);
            end
            MAX: begin
                result = (input1 > input2) ? input1 : input2;
            end
            MIN: begin
                result = (input1 < input2) ? input1 : input2;
            end
            ADD: begin
                result = input1 + input2;
                overflow = (input1[7] == input2[7]) && (result[7] != input1[7]);
            end
            SLL: begin
                result = input1 << shiftValue;
            end
            SUB: begin
                result = input1 - input2;
                overflow = (input1[7] != input2[7]) && (result[7] != input1[7]);
            end
            XOR: begin
                result = input1 ^ input2;
            end
            XNOR: begin
                result = ~(input1 ^ input2);
            end
            SRA: begin
                result = $signed(input1) >>> shiftValue;
            end
            default: result = 8'b0;
        endcase
        zeroFlag = (result == 8'b0);
        signFlag = result[7];
    end

endmodule