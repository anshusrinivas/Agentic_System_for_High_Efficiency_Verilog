`timescale 1ns / 1ps

// Generated ALU Module
// Style: FUNCTION
// Bit width: 8
// Operations: ROL, ROR, MAX, MIN, SRL, PASSB, AND
// Flags: carry, zero, overflow

module ALU_1579W8_b60d197f(
    input  wire [3:0]  opcode,
    input  wire [7:0] input1,
    input  wire [7:0] input2,
    input  wire [4:0]       shiftValue,
    output wire [7:0] result
    ,output wire carryFlag
    ,output wire zeroFlag
    ,output wire overFlowFlag
);

    function [7:0] rol;
        input [7:0] a;
        input [4:0] sh;
        begin
            rol = (a << sh) | (a >> (8-sh));
        end
    endfunction

    function [7:0] ror;
        input [7:0] a;
        input [4:0] sh;
        begin
            ror = (a >> sh) | (a << (8-sh));
        end
    endfunction

    // Operation codes
    localparam ROL = 4'd0;
    localparam ROR = 4'd1;
    localparam MAX = 4'd2;
    localparam MIN = 4'd3;
    localparam SRL = 4'd4;
    localparam PASSB = 4'd5;
    localparam AND = 4'd6;

    // Combinational logic
    always @(*) begin
        case (opcode)
            ROL: begin
                result = rol(input1, shiftValue);
            end
            ROR: begin
                result = ror(input1, shiftValue);
            end
            MAX: begin
                result = (input1 > input2) ? input1 : input2;
            end
            MIN: begin
                result = (input1 < input2) ? input1 : input2;
            end
            SRL: begin
                result = input1 >> shiftValue;
            end
            PASSB: begin
                result = input2;
            end
            AND: begin
                result = input1 & input2;
            end
            default: result = 8'b0;
        endcase
        zeroFlag = (result == 8'b0);
    end

endmodule