`timescale 1ns / 1ps

// Generated ALU Module
// Style: MODULAR
// Bit width: 128
// Operations: SLL, MIN, PASSB, XNOR, SNE, DIV, SGE, ADD, ROL, NAND, SRA, SUB
// Flags: carry, zero, overflow, sign

module ALU_1842W128_b3f6b71c(
    input  wire [3:0]  opcode,
    input  wire [127:0] input1,
    input  wire [127:0] input2,
    input  wire [4:0]       shiftValue,
    output reg  [127:0] result
    ,output reg  carryFlag
    ,output reg  zeroFlag
    ,output reg  overFlowFlag
    ,output reg  signFlag
);

    // Operation codes
    localparam SLL = 4'd0;
    localparam MIN = 4'd1;
    localparam PASSB = 4'd2;
    localparam XNOR = 4'd3;
    localparam SNE = 4'd4;
    localparam DIV = 4'd5;
    localparam SGE = 4'd6;
    localparam ADD = 4'd7;
    localparam ROL = 4'd8;
    localparam NAND = 4'd9;
    localparam SRA = 4'd10;
    localparam SUB = 4'd11;

    // Combinational logic
    always @(*) begin
        case (opcode)
            SLL: begin
                result = input1 << shiftValue;
            end
            MIN: begin
                result = (input1 < input2) ? input1 : input2;
            end
            PASSB: begin
                result = input2;
            end
            XNOR: begin
                result = ~(input1 ^ input2);
            end
            SNE: begin
            end
            DIV: begin
                result = (input2 != 0) ? input1 / input2 : 128'b0;
            end
            SGE: begin
            end
            ADD: begin
                result = input1 + input2;
                overflow = (input1[127] == input2[127]) && (result[127] != input1[127]);
            end
            ROL: begin
                result = rol(input1, shiftValue);
            end
            NAND: begin
                result = ~(input1 & input2);
            end
            SRA: begin
                result = $signed(input1) >>> shiftValue;
            end
            SUB: begin
                result = input1 - input2;
                overflow = (input1[127] != input2[127]) && (result[127] != input1[127]);
            end
            default: result = 128'b0;
        endcase
        zeroFlag = (result == 128'b0);
        signFlag = result[127];
    end

endmodule