`timescale 1ns / 1ps

// Generated ALU Module
// Style: FUNCTION
// Bit width: 128
// Operations: ROL, ROR, MAX, MIN
// Flags: carry, zero, overflow

module ALU_0807W128_466836be(
    input  wire [3:0]  opcode,
    input  wire [127:0] input1,
    input  wire [127:0] input2,
    input  wire [4:0]       shiftValue,
    output wire [127:0] result
    ,output wire carryFlag
    ,output wire zeroFlag
    ,output wire overFlowFlag
);

    function [127:0] rol;
        input [127:0] a;
        input [4:0] sh;
        begin
            rol = (a << sh) | (a >> (128-sh));
        end
    endfunction

    function [127:0] ror;
        input [127:0] a;
        input [4:0] sh;
        begin
            ror = (a >> sh) | (a << (128-sh));
        end
    endfunction

    // Operation codes
    localparam ROL = 4'd0;
    localparam ROR = 4'd1;
    localparam MAX = 4'd2;
    localparam MIN = 4'd3;

    // Combinational logic
    always @(*) begin
        case (opcode)
            ROL: begin
                result = rol(input1, shiftValue);
            end
            ROR: begin
                result = ror(input1, shiftValue);
            end
            MAX: begin
                result = (input1 > input2) ? input1 : input2;
            end
            MIN: begin
                result = (input1 < input2) ? input1 : input2;
            end
            default: result = 128'b0;
        endcase
        zeroFlag = (result == 128'b0);
    end

endmodule