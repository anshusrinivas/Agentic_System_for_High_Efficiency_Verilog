`timescale 1ns / 1ps

// Generated ALU Module
// Style: MODULAR
// Bit width: 64
// Operations: AND, MUL, SLTU, NOR, DIV, SRA, ROR, XNOR, SGT, XOR, ADD, SUB, SLT, SEQ
// Flags: carry, zero, overflow, sign

module ALU_1768W64_44f23a52(
    input  wire [3:0]  opcode,
    input  wire [63:0] input1,
    input  wire [63:0] input2,
    input  wire [4:0]       shiftValue,
    output reg  [63:0] result
    ,output reg  carryFlag
    ,output reg  zeroFlag
    ,output reg  overFlowFlag
    ,output reg  signFlag
);

    // Operation codes
    localparam AND = 4'd0;
    localparam MUL = 4'd1;
    localparam SLTU = 4'd2;
    localparam NOR = 4'd3;
    localparam DIV = 4'd4;
    localparam SRA = 4'd5;
    localparam ROR = 4'd6;
    localparam XNOR = 4'd7;
    localparam SGT = 4'd8;
    localparam XOR = 4'd9;
    localparam ADD = 4'd10;
    localparam SUB = 4'd11;
    localparam SLT = 4'd12;
    localparam SEQ = 4'd13;

    // Combinational logic
    always @(*) begin
        case (opcode)
            AND: begin
                result = input1 & input2;
            end
            MUL: begin
                result = input1 * input2;
            end
            SLTU: begin
            end
            NOR: begin
                result = ~(input1 | input2);
            end
            DIV: begin
                result = (input2 != 0) ? input1 / input2 : 64'b0;
            end
            SRA: begin
                result = $signed(input1) >>> shiftValue;
            end
            ROR: begin
                result = ror(input1, shiftValue);
            end
            XNOR: begin
                result = ~(input1 ^ input2);
            end
            SGT: begin
            end
            XOR: begin
                result = input1 ^ input2;
            end
            ADD: begin
                result = input1 + input2;
                overflow = (input1[63] == input2[63]) && (result[63] != input1[63]);
            end
            SUB: begin
                result = input1 - input2;
                overflow = (input1[63] != input2[63]) && (result[63] != input1[63]);
            end
            SLT: begin
            end
            SEQ: begin
            end
            default: result = 64'b0;
        endcase
        zeroFlag = (result == 64'b0);
        signFlag = result[63];
    end

endmodule