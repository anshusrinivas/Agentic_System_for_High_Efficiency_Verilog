`timescale 1ns / 1ps

// Generated ALU Module
// Style: OPTIMIZED
// Bit width: 64
// Operations: ADD, SUB, AND, OR, SLL, NOR, ROL, SRL, SRA
// Flags: carry, zero, sign

module ALU_1892W64_8aee8688(
    input  wire [3:0]  opcode,
    input  wire [63:0] input1,
    input  wire [63:0] input2,
    input  wire [4:0]       shiftValue,
    output reg  [63:0] result
    ,output reg  carryFlag
    ,output reg  zeroFlag
    ,output reg  signFlag
);

    // Operation codes
    localparam ADD = 4'd0;
    localparam SUB = 4'd1;
    localparam AND = 4'd2;
    localparam OR = 4'd3;
    localparam SLL = 4'd4;
    localparam NOR = 4'd5;
    localparam ROL = 4'd6;
    localparam SRL = 4'd7;
    localparam SRA = 4'd8;

    // Internal signals
    wire [64:0] sum = (opcode == SUB) ? 
                             {1'b0, input1} - {1'b0, input2} : 
                             {1'b0, input1} + {1'b0, input2};

    // Combinational logic
    always @(*) begin
        case (opcode)
            ADD: begin
                result = input1 + input2;
                
            end
            SUB: begin
                result = input1 - input2;
                
            end
            AND: begin
                result = input1 & input2;
            end
            OR: begin
                result = input1 | input2;
            end
            SLL: begin
                result = input1 << shiftValue;
            end
            NOR: begin
                result = ~(input1 | input2);
            end
            ROL: begin
                result = rol(input1, shiftValue);
            end
            SRL: begin
                result = input1 >> shiftValue;
            end
            SRA: begin
                result = $signed(input1) >>> shiftValue;
            end
            default: result = 64'b0;
        endcase
        zeroFlag = (result == 64'b0);
        signFlag = result[63];
    end

endmodule