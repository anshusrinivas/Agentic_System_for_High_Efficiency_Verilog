`timescale 1ns / 1ps

// Generated ALU Module
// Style: STANDARD
// Bit width: 64
// Operations: ADD, SUB, AND, OR, NAND, ROL, MUL, DIV, MIN, MAX
// Flags: carry, zero, overflow, sign

module ALU_1305W64_efa3d54a(
    input  wire [3:0]  opcode,
    input  wire [63:0] input1,
    input  wire [63:0] input2,
    input  wire [4:0]       shiftValue,
    output wire [63:0] result
    ,output wire carryFlag
    ,output wire zeroFlag
    ,output wire overFlowFlag
    ,output wire signFlag
);

    // Operation codes
    localparam ADD = 4'd0;
    localparam SUB = 4'd1;
    localparam AND = 4'd2;
    localparam OR = 4'd3;
    localparam NAND = 4'd4;
    localparam ROL = 4'd5;
    localparam MUL = 4'd6;
    localparam DIV = 4'd7;
    localparam MIN = 4'd8;
    localparam MAX = 4'd9;

    // Internal signals
    wire [64:0] sum = (opcode == SUB) ? 
                             {1'b0, input1} - {1'b0, input2} : 
                             {1'b0, input1} + {1'b0, input2};

    // Combinational logic
    always @(*) begin
        case (opcode)
            ADD: begin
                result = input1 + input2;
                overflow = (input1[63] == input2[63]) && (result[63] != input1[63]);
            end
            SUB: begin
                result = input1 - input2;
                overflow = (input1[63] != input2[63]) && (result[63] != input1[63]);
            end
            AND: begin
                result = input1 & input2;
            end
            OR: begin
                result = input1 | input2;
            end
            NAND: begin
                result = ~(input1 & input2);
            end
            ROL: begin
                result = rol(input1, shiftValue);
            end
            MUL: begin
                result = input1 * input2;
            end
            DIV: begin
                result = (input2 != 0) ? input1 / input2 : 64'b0;
            end
            MIN: begin
                result = (input1 < input2) ? input1 : input2;
            end
            MAX: begin
                result = (input1 > input2) ? input1 : input2;
            end
            default: result = 64'b0;
        endcase
        zeroFlag = (result == 64'b0);
        signFlag = result[63];
    end

endmodule