`timescale 1ns / 1ps

// Generated ALU Module
// Style: STANDARD
// Bit width: 8
// Operations: ADD, SUB, AND, OR, MUL, MAX, NOR, SRA, DIV
// Flags: carry

module ALU_0611W8_72ce2b97(
    input  wire [3:0]  opcode,
    input  wire [7:0] input1,
    input  wire [7:0] input2,
    input  wire [4:0]       shiftValue,
    output wire [7:0] result
    ,output wire carryFlag
);

    // Operation codes
    localparam ADD = 4'd0;
    localparam SUB = 4'd1;
    localparam AND = 4'd2;
    localparam OR = 4'd3;
    localparam MUL = 4'd4;
    localparam MAX = 4'd5;
    localparam NOR = 4'd6;
    localparam SRA = 4'd7;
    localparam DIV = 4'd8;

    // Internal signals
    wire [8:0] sum = (opcode == SUB) ? 
                             {1'b0, input1} - {1'b0, input2} : 
                             {1'b0, input1} + {1'b0, input2};

    // Combinational logic
    always @(*) begin
        case (opcode)
            ADD: begin
                result = input1 + input2;
                
            end
            SUB: begin
                result = input1 - input2;
                
            end
            AND: begin
                result = input1 & input2;
            end
            OR: begin
                result = input1 | input2;
            end
            MUL: begin
                result = input1 * input2;
            end
            MAX: begin
                result = (input1 > input2) ? input1 : input2;
            end
            NOR: begin
                result = ~(input1 | input2);
            end
            SRA: begin
                result = $signed(input1) >>> shiftValue;
            end
            DIV: begin
                result = (input2 != 0) ? input1 / input2 : 8'b0;
            end
            default: result = 8'b0;
        endcase
    end

endmodule