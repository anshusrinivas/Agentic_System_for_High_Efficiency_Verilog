`timescale 1ns / 1ps

// Generated ALU Module
// Style: MODULAR
// Bit width: 128
// Operations: NAND, ROR, ROL, MAX, PASSB, SLL, NOR, SNE, SRA, ADD, AND
// Flags: carry, zero, overflow

module ALU_0360W128_6ee44902(
    input  wire [3:0]  opcode,
    input  wire [127:0] input1,
    input  wire [127:0] input2,
    input  wire [4:0]       shiftValue,
    output reg  [127:0] result
    ,output reg  carryFlag
    ,output reg  zeroFlag
    ,output reg  overFlowFlag
);

    // Operation codes
    localparam NAND = 4'd0;
    localparam ROR = 4'd1;
    localparam ROL = 4'd2;
    localparam MAX = 4'd3;
    localparam PASSB = 4'd4;
    localparam SLL = 4'd5;
    localparam NOR = 4'd6;
    localparam SNE = 4'd7;
    localparam SRA = 4'd8;
    localparam ADD = 4'd9;
    localparam AND = 4'd10;

    // Combinational logic
    always @(*) begin
        case (opcode)
            NAND: begin
                result = ~(input1 & input2);
            end
            ROR: begin
                result = ror(input1, shiftValue);
            end
            ROL: begin
                result = rol(input1, shiftValue);
            end
            MAX: begin
                result = (input1 > input2) ? input1 : input2;
            end
            PASSB: begin
                result = input2;
            end
            SLL: begin
                result = input1 << shiftValue;
            end
            NOR: begin
                result = ~(input1 | input2);
            end
            SNE: begin
            end
            SRA: begin
                result = $signed(input1) >>> shiftValue;
            end
            ADD: begin
                result = input1 + input2;
                overflow = (input1[127] == input2[127]) && (result[127] != input1[127]);
            end
            AND: begin
                result = input1 & input2;
            end
            default: result = 128'b0;
        endcase
        zeroFlag = (result == 128'b0);
    end

endmodule