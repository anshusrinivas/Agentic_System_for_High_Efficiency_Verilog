`timescale 1ns / 1ps

// Generated ALU Module
// Style: MODULAR
// Bit width: 128
// Operations: SRL, XNOR, ROR, SLL, OR, SUB, SGT, MAX, NAND, ADD, MIN
// Flags: carry, zero, overflow, sign

module ALU_0344W128_9bdb9ae1(
    input  wire [3:0]  opcode,
    input  wire [127:0] input1,
    input  wire [127:0] input2,
    input  wire [4:0]       shiftValue,
    output reg  [127:0] result
    ,output reg  carryFlag
    ,output reg  zeroFlag
    ,output reg  overFlowFlag
    ,output reg  signFlag
);

    // Operation codes
    localparam SRL = 4'd0;
    localparam XNOR = 4'd1;
    localparam ROR = 4'd2;
    localparam SLL = 4'd3;
    localparam OR = 4'd4;
    localparam SUB = 4'd5;
    localparam SGT = 4'd6;
    localparam MAX = 4'd7;
    localparam NAND = 4'd8;
    localparam ADD = 4'd9;
    localparam MIN = 4'd10;

    // Combinational logic
    always @(*) begin
        case (opcode)
            SRL: begin
                result = input1 >> shiftValue;
            end
            XNOR: begin
                result = ~(input1 ^ input2);
            end
            ROR: begin
                result = ror(input1, shiftValue);
            end
            SLL: begin
                result = input1 << shiftValue;
            end
            OR: begin
                result = input1 | input2;
            end
            SUB: begin
                result = input1 - input2;
                overflow = (input1[127] != input2[127]) && (result[127] != input1[127]);
            end
            SGT: begin
            end
            MAX: begin
                result = (input1 > input2) ? input1 : input2;
            end
            NAND: begin
                result = ~(input1 & input2);
            end
            ADD: begin
                result = input1 + input2;
                overflow = (input1[127] == input2[127]) && (result[127] != input1[127]);
            end
            MIN: begin
                result = (input1 < input2) ? input1 : input2;
            end
            default: result = 128'b0;
        endcase
        zeroFlag = (result == 128'b0);
        signFlag = result[127];
    end

endmodule